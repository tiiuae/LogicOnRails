module module_eg #(

)(
    input  logic       i_clk,
    input  logic       i_rst_n
);

////////////////////////////////////////
//                signals
////////////////////////////////////////

////////////////////////////////////////
//                <name>
////////////////////////////////////////

always_ff @(posedge i_clk or negedge i_rst_n)
begin
    if(i_rst_n == 1'b0) begin
    end else begin
    end
end

always_comb 
begin
end

////////////////////////////////////////
//                outputs
////////////////////////////////////////

endmodule
