package iface_tb_pkg;

    localparam AVALON_ST_BUS_WIDTH = 32;

    localparam AXI_ST_BUS_WIDTH    = 96;
    localparam AXI_ST_USR_WIDTH    = 16;

    localparam AXI4_ADDR_WIDTH    = 16;
    localparam AXI4_DATA_WIDTH    = 32;
    localparam AXI4_WRBURST_VAL   = 1;
    localparam AXI4_WRLEN_VAL     = 7;
    localparam AXI4_WRPROT_VAL    = 0;
    localparam AXI4_ADDR_RND      = 0;

endpackage
