`timescale 1ns/1ps

module pll_2 (
    input  logic       refclk,
    output logic       locked,
    input  logic       rst,
    output logic       outclk_0
);


endmodule
