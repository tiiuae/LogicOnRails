`timescale 1ns/1ps  
package io_pkg;


endpackage
